function incremnt_gcm (input [127:0] j0);
	begin 
		incremnt_gcm = j0 + 1 ; 
	end
endfunction : 