module tb_aes_sbox ();

/**********************************************************************
* Inputs as registers
**********************************************************************/
	reg [31:0] i_wrd_sbox;

/**********************************************************************
* output as wires
**********************************************************************/
	wire [31:0] o_wrd_sbox;

/**********************************************************************
* DUT instantiation
**********************************************************************/

	aes_sbox DUT (
		.i_wrd_sbox(i_wrd_sbox),
		.o_wrd_sbox(o_wrd_sbox)
	);
/**********************************************************************
* Stimulus here
**********************************************************************/

	initial
		begin
			repeat (5)
				begin
					i_wrd_sbox = $random();
					#5;
				end
		end
endmodule