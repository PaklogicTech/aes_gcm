module tb_aes_inv_sbox ();

/**********************************************************************
* Inputs as registers 
**********************************************************************/
reg  [31 : 0] i_inv_wrd_sbox; 

/**********************************************************************
* output as wires 
**********************************************************************/
wire [31 : 0] o_inv_wrd_sbox; 

/**********************************************************************
* DUT instantiation 
**********************************************************************/

aes_inv_sbox DUT(

                   .i_inv_wrd_sbox(i_inv_wrd_sbox),
                   .o_inv_wrd_sbox(o_inv_wrd_sbox)
                   );
/**********************************************************************
* Stimulus here
**********************************************************************/

initial
begin 
	i_inv_wrd_sbox = $random();
end
endmodule