module tb_mul_128_module ();


/**********************************************************************
* Inputs as register
**********************************************************************/

	reg [127:0] B;
	reg [127:0] A;

/**********************************************************************
* outputs as wire
**********************************************************************/

	wire [255:0] mul_128;

	mul_128_module DUT(
		.B(B),
		.A(A),
		.mul_128(mul_128)
	);


	task run_sim();
		begin
			A='d10;
			B='d20;
//			A=$random();
//			B=$random();
		end
	endtask : run_sim

	initial 
	begin 
		run_sim();
	end

endmodule